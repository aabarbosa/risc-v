module vJTAG_interface (
	input logic [7:0] r [0:31]
);


endmodule

